V2 VDD GND DC 12
.end
